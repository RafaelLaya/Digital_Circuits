/*	ROM module that stores Sprite for fireball
 *		Outputs:
 *			fireball_sprite		- Sprite for fireball
 *
 * Position [x][y][{r,g,b}] contains pixel at (x, y) where r, g, b are 8 bits each
 * (0, 0) is at the top-left
 * Width 45, Height 36, Color-depth 24
*/

module ROM_fireball_sprite (fireball_sprite);
	output logic [35:0][23:0] fireball_sprite [44:0];

	assign fireball_sprite[0] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[1] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[2] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[3] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[4] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[5] =  { 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[6] =  { 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[7] =  { 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0 };
	assign fireball_sprite[8] =  { 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0 };
	assign fireball_sprite[9] =  { 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd0, 24'd0 };
	assign fireball_sprite[10] =  { 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd0, 24'd0 };
	assign fireball_sprite[11] =  { 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd0, 24'd0 };
	assign fireball_sprite[12] =  { 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16777215, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd0, 24'd0 };
	assign fireball_sprite[13] =  { 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd0, 24'd0 };
	assign fireball_sprite[14] =  { 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd0, 24'd0 };
	assign fireball_sprite[15] =  { 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd0, 24'd0 };
	assign fireball_sprite[16] =  { 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd0, 24'd0 };
	assign fireball_sprite[17] =  { 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd0, 24'd0 };
	assign fireball_sprite[18] =  { 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd0, 24'd0 };
	assign fireball_sprite[19] =  { 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd0, 24'd0 };
	assign fireball_sprite[20] =  { 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd0, 24'd0 };
	assign fireball_sprite[21] =  { 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0 };
	assign fireball_sprite[22] =  { 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[23] =  { 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16772096, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[24] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[25] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[26] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[27] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[28] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[29] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[30] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[31] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[32] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[33] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd6356992, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[34] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[35] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[36] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16743424, 24'd16743424, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[37] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[38] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[39] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[40] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[41] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[42] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[43] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign fireball_sprite[44] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };

endmodule // ROM_fireball_sprite