/*	ROM module that stores Sprite for the floor
 *		Outputs:
 *			floor_sprite		- Sprite for the floor
 *
 * Position [x][y][{r,g,b}] contains pixel at (x, y) where r, g, b are 8 bits each
 * (0, 0) is at the top-left
 * Width 640, Height 8, Color-depth 24
*/
module ROM_floor_sprite(floor_sprite);
	output logic [7:0][23:0] floor_sprite [639:0];

	assign floor_sprite[0] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[1] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[2] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[3] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[4] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[5] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[6] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[7] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[8] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[9] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[10] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[11] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[12] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[13] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[14] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[15] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[16] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[17] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[18] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[19] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[20] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[21] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[22] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[23] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[24] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[25] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[26] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[27] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[28] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[29] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[30] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[31] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[32] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[33] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[34] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[35] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[36] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[37] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[38] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[39] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[40] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[41] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[42] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[43] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[44] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[45] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[46] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[47] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[48] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[49] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[50] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[51] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[52] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[53] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[54] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[55] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[56] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[57] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[58] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[59] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[60] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[61] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[62] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[63] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[64] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[65] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[66] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[67] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[68] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[69] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[70] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[71] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[72] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[73] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[74] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[75] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[76] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[77] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[78] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[79] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[80] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[81] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[82] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[83] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[84] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[85] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[86] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[87] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[88] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[89] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[90] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[91] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[92] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[93] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[94] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[95] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[96] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[97] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[98] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[99] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[100] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[101] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[102] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[103] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[104] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[105] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[106] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[107] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[108] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[109] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[110] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[111] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[112] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[113] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[114] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[115] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[116] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[117] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[118] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[119] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[120] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[121] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[122] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[123] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[124] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[125] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[126] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[127] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[128] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[129] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[130] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[131] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[132] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[133] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[134] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[135] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[136] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[137] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[138] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[139] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[140] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[141] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[142] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[143] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[144] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[145] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[146] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[147] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[148] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[149] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[150] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[151] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[152] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[153] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[154] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[155] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[156] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[157] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[158] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[159] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[160] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[161] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[162] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[163] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[164] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[165] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[166] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[167] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[168] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[169] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[170] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[171] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[172] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[173] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[174] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[175] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[176] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[177] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[178] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[179] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[180] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[181] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[182] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[183] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[184] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[185] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[186] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[187] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[188] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[189] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[190] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[191] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[192] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[193] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[194] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[195] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[196] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[197] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[198] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[199] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[200] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[201] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[202] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[203] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[204] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[205] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[206] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[207] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[208] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[209] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[210] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[211] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[212] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[213] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[214] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[215] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[216] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[217] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[218] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[219] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[220] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[221] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[222] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[223] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[224] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[225] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[226] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[227] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[228] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[229] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[230] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[231] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[232] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[233] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[234] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[235] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[236] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[237] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[238] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[239] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[240] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[241] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[242] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[243] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[244] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[245] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[246] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[247] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[248] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[249] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[250] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[251] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[252] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[253] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[254] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[255] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[256] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[257] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[258] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[259] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[260] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[261] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[262] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[263] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[264] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[265] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[266] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[267] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[268] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[269] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[270] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[271] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[272] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[273] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[274] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[275] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[276] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[277] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[278] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[279] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[280] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[281] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[282] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[283] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[284] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[285] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[286] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[287] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[288] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[289] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[290] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[291] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[292] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[293] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[294] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[295] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[296] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[297] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[298] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[299] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[300] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[301] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[302] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[303] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[304] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[305] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[306] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[307] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[308] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[309] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[310] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[311] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[312] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[313] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[314] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[315] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[316] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[317] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[318] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[319] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[320] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[321] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[322] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[323] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[324] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[325] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[326] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[327] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[328] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[329] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[330] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[331] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[332] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[333] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[334] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[335] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[336] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[337] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[338] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[339] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[340] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[341] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[342] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[343] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[344] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[345] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[346] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[347] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[348] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[349] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[350] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[351] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[352] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[353] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[354] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[355] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[356] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[357] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[358] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[359] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[360] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[361] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[362] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[363] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[364] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[365] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[366] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[367] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[368] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[369] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[370] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[371] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[372] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[373] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[374] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[375] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[376] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[377] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[378] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[379] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[380] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[381] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[382] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[383] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[384] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[385] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[386] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[387] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[388] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[389] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[390] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[391] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[392] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[393] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[394] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[395] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[396] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[397] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[398] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[399] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[400] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[401] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[402] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[403] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[404] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[405] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[406] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[407] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[408] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[409] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[410] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[411] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[412] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[413] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[414] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[415] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[416] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[417] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[418] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[419] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[420] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[421] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[422] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[423] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[424] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[425] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[426] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[427] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[428] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[429] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[430] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[431] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[432] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[433] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[434] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[435] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[436] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[437] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[438] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[439] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[440] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[441] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[442] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[443] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[444] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[445] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[446] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[447] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[448] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[449] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[450] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[451] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[452] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[453] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[454] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[455] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[456] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[457] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[458] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[459] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[460] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[461] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[462] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[463] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[464] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[465] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[466] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[467] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[468] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[469] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[470] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[471] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[472] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[473] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[474] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[475] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[476] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[477] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[478] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[479] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[480] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[481] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[482] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[483] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[484] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[485] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[486] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[487] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[488] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[489] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[490] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[491] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[492] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[493] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[494] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[495] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[496] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[497] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[498] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[499] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[500] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[501] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[502] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[503] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[504] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[505] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[506] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[507] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[508] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[509] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[510] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[511] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[512] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[513] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[514] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[515] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[516] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[517] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[518] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[519] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[520] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[521] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[522] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[523] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[524] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[525] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[526] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[527] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[528] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[529] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[530] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[531] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[532] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[533] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[534] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[535] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[536] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[537] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[538] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[539] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[540] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[541] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[542] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[543] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[544] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[545] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[546] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[547] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[548] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[549] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[550] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[551] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[552] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[553] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[554] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[555] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[556] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[557] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[558] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[559] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[560] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[561] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[562] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[563] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[564] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[565] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[566] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[567] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[568] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[569] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[570] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[571] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[572] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[573] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[574] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[575] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[576] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[577] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[578] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[579] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[580] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[581] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[582] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[583] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[584] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[585] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[586] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[587] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[588] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[589] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[590] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[591] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[592] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[593] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[594] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[595] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[596] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[597] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[598] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[599] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[600] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[601] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[602] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[603] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[604] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[605] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[606] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[607] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[608] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[609] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[610] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[611] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[612] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[613] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[614] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[615] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280 };
	assign floor_sprite[616] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[617] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[618] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[619] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[620] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0 };
	assign floor_sprite[621] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[622] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[623] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[624] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[625] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[626] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[627] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[628] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[629] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[630] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[631] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[632] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[633] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[634] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[635] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[636] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[637] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0, 24'd0, 24'd0 };
	assign floor_sprite[638] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
	assign floor_sprite[639] =  { 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd6324280, 24'd0 };
		
endmodule // ROM_floor_sprite