/*	ROM module that stores Sprite #1 for dyno in running position
 *		Outputs:
 *			dyno_running_sprite1			- sprite #1 for dyno in running position
 *
 * Position [x][y][{r,g,b}] contains pixel at (x, y) where r, g, b are 8 bits each
 * (0, 0) is at the top-left
 * Width 32, Height 32, Color-depth 24
*/
module ROM_dyno_running_sprite1(dyno_running_sprite1);

	output logic [31:0][23:0] dyno_running_sprite1 [0:31];
		
	assign dyno_running_sprite1[0] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_running_sprite1[1] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_running_sprite1[2] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_running_sprite1[3] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd0 };
	assign dyno_running_sprite1[4] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd0 };
	assign dyno_running_sprite1[5] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd0 };
	assign dyno_running_sprite1[6] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680 };
	assign dyno_running_sprite1[7] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680 };
	assign dyno_running_sprite1[8] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680 };
	assign dyno_running_sprite1[9] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite1[10] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite1[11] =  { 24'd8323072, 24'd8323072, 24'd8323072, 24'd8323072, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite1[12] =  { 24'd8323072, 24'd8323072, 24'd8323072, 24'd8323072, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite1[13] =  { 24'd8323072, 24'd8323072, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd10526880, 24'd10526880, 24'd10526880, 24'd5011456, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite1[14] =  { 24'd8323072, 24'd8323072, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite1[15] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite1[16] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite1[17] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite1[18] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd8323072, 24'd8323072, 24'd8323072, 24'd8323072, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd16757375, 24'd16757375, 24'd16711680, 24'd16711680, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite1[19] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd8323072, 24'd8323072, 24'd8323072, 24'd8323072, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd16757375, 24'd16757375, 24'd16711680, 24'd16711680, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite1[20] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd8323072, 24'd8323072, 24'd0, 24'd0, 24'd0, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16757375, 24'd16757375, 24'd38143, 24'd38143, 24'd16757375, 24'd5011456, 24'd0, 24'd0 };
	assign dyno_running_sprite1[21] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd8323072, 24'd8323072, 24'd0, 24'd0, 24'd0, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16757375, 24'd16757375, 24'd38143, 24'd38143, 24'd16757375, 24'd5011456, 24'd0, 24'd0 };
	assign dyno_running_sprite1[22] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd8323072, 24'd8323072, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16757375, 24'd16757375, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_running_sprite1[23] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16757375, 24'd16757375, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_running_sprite1[24] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16757375, 24'd16757375, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_running_sprite1[25] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16757375, 24'd16757375, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_running_sprite1[26] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16757375, 24'd16757375, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_running_sprite1[27] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd16711680, 24'd16711680, 24'd0, 24'd0 };
	assign dyno_running_sprite1[28] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0 };
	assign dyno_running_sprite1[29] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_running_sprite1[30] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_running_sprite1[31] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
		
endmodule // ROM_dyno_running_sprite1