/*	ROM module that stores Sprite #0 for dyno in ducking position
 *		Outputs:
 *			dyno_ducking0_sprite			- sprite #0 for dyno in ducking position
 *
 * Position [x][y][{r,g,b}] contains pixel at (x, y) where r, g, b are 8 bits each
 * (0, 0) is at the top-left
 * Width 32, Height 32, Color-depth 24
*/

module ROM_dyno_ducking0_sprite(dyno_ducking0_sprite);
	output logic [31:0][23:0] dyno_ducking0_sprite [0:31];

		
	assign dyno_ducking0_sprite[0] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[1] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[2] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[3] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[4] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[5] =  { 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[6] =  { 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[7] =  { 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[8] =  { 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[9] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[10] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[11] =  { 24'd8323072, 24'd8323072, 24'd8323072, 24'd16757375, 24'd16757375, 24'd5011456, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[12] =  { 24'd8323072, 24'd8323072, 24'd8323072, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd10526880, 24'd10526880, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[13] =  { 24'd8323072, 24'd8323072, 24'd0, 24'd0, 24'd0, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[14] =  { 24'd8323072, 24'd8323072, 24'd0, 24'd0, 24'd0, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[15] =  { 24'd8323072, 24'd8323072, 24'd0, 24'd0, 24'd0, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[16] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[17] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[18] =  { 24'd0, 24'd0, 24'd0, 24'd8323072, 24'd8323072, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd16757375, 24'd16711680, 24'd16711680, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[19] =  { 24'd0, 24'd0, 24'd0, 24'd8323072, 24'd8323072, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd16757375, 24'd16711680, 24'd16711680, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[20] =  { 24'd0, 24'd0, 24'd0, 24'd8323072, 24'd8323072, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd0, 24'd16711680, 24'd16711680, 24'd16757375, 24'd16757375, 24'd38143, 24'd38143, 24'd5011456, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[21] =  { 24'd0, 24'd0, 24'd0, 24'd8323072, 24'd8323072, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd0, 24'd16711680, 24'd16711680, 24'd16757375, 24'd16757375, 24'd38143, 24'd38143, 24'd5011456, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[22] =  { 24'd0, 24'd0, 24'd0, 24'd8323072, 24'd8323072, 24'd0, 24'd16757375, 24'd16757375, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[23] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16757375, 24'd16757375, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[24] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16757375, 24'd16757375, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[25] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16757375, 24'd16757375, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[26] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[27] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[28] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[29] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[30] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_ducking0_sprite[31] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };

endmodule // ROM_dyno_ducking0_sprite