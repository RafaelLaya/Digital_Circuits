/*	ROM module that stores Sprite #0 for witch
 *		Outputs:
 *			witch_sprite0		- Sprite #0 for witch
 *
 * Position [x][y][{r,g,b}] contains pixel at (x, y) where r, g, b are 8 bits each
 * (0, 0) is at the top-left
 * Width 45, Height 36, Color-depth 24
*/

module ROM_witch_sprite0(witch_sprite0);

	output logic [35:0][23:0] witch_sprite0[44:0];

	assign witch_sprite0[0] =  { 24'd0, 24'd0, 24'd0, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[1] =  { 24'd0, 24'd0, 24'd0, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[2] =  { 24'd0, 24'd0, 24'd0, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[3] =  { 24'd0, 24'd0, 24'd0, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[4] =  { 24'd0, 24'd0, 24'd0, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[5] =  { 24'd0, 24'd0, 24'd0, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[6] =  { 24'd0, 24'd0, 24'd0, 24'd6438947, 24'd6438947, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[7] =  { 24'd0, 24'd0, 24'd0, 24'd6438947, 24'd6438947, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[8] =  { 24'd0, 24'd0, 24'd0, 24'd6438947, 24'd6438947, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[9] =  { 24'd0, 24'd0, 24'd0, 24'd6438947, 24'd6438947, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[10] =  { 24'd0, 24'd0, 24'd0, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd16777215, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd16711680, 24'd16711680, 24'd16711680, 24'd5291375, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[11] =  { 24'd0, 24'd0, 24'd0, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd6438947, 24'd16777215, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd16711680, 24'd16711680, 24'd16711680, 24'd5291375, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[12] =  { 24'd0, 24'd0, 24'd0, 24'd6438947, 24'd6438947, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd16711680, 24'd16711680, 24'd5291375, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[13] =  { 24'd0, 24'd0, 24'd0, 24'd6438947, 24'd6438947, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd16777215, 24'd16777215, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[14] =  { 24'd0, 24'd0, 24'd0, 24'd6438947, 24'd6438947, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd16777215, 24'd16777215, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[15] =  { 24'd0, 24'd0, 24'd0, 24'd6438947, 24'd6438947, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd16777215, 24'd16777215, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd9607588, 24'd9607588, 24'd9607588, 24'd1118481, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[16] =  { 24'd0, 24'd0, 24'd0, 24'd6438947, 24'd6438947, 24'd6438947, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[17] =  { 24'd0, 24'd0, 24'd0, 24'd6438947, 24'd6438947, 24'd6438947, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[18] =  { 24'd0, 24'd0, 24'd0, 24'd6438947, 24'd6438947, 24'd6438947, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[19] =  { 24'd0, 24'd0, 24'd0, 24'd6438947, 24'd6438947, 24'd4564320, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[20] =  { 24'd0, 24'd0, 24'd0, 24'd6438947, 24'd6438947, 24'd4564320, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[21] =  { 24'd0, 24'd0, 24'd0, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd5291375, 24'd5291375, 24'd5291375, 24'd5291375, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd9607588, 24'd9607588, 24'd9607588, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0 };
	assign witch_sprite0[22] =  { 24'd0, 24'd0, 24'd0, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd3092270, 24'd3092270, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784 };
	assign witch_sprite0[23] =  { 24'd0, 24'd0, 24'd0, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4564320, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd3092270, 24'd3092270, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784 };
	assign witch_sprite0[24] =  { 24'd0, 24'd0, 24'd0, 24'd4564320, 24'd4564320, 24'd4564320, 24'd6438947, 24'd6438947, 24'd6438947, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784 };
	assign witch_sprite0[25] =  { 24'd0, 24'd0, 24'd0, 24'd4564320, 24'd4564320, 24'd4564320, 24'd6438947, 24'd6438947, 24'd6438947, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784 };
	assign witch_sprite0[26] =  { 24'd0, 24'd0, 24'd0, 24'd4564320, 24'd4564320, 24'd4564320, 24'd6438947, 24'd6438947, 24'd6438947, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784 };
	assign witch_sprite0[27] =  { 24'd0, 24'd0, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd4402784, 24'd4402784, 24'd4402784, 24'd3745617, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784 };
	assign witch_sprite0[28] =  { 24'd0, 24'd0, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784 };
	assign witch_sprite0[29] =  { 24'd0, 24'd0, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd9607588, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784 };
	assign witch_sprite0[30] =  { 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9607588, 24'd9607588, 24'd9607588, 24'd0, 24'd0, 24'd3745617, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0 };
	assign witch_sprite0[31] =  { 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[32] =  { 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[33] =  { 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[34] =  { 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[35] =  { 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[36] =  { 24'd0, 24'd0, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[37] =  { 24'd0, 24'd0, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[38] =  { 24'd0, 24'd0, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd4402784, 24'd4402784, 24'd4402784, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[39] =  { 24'd0, 24'd0, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[40] =  { 24'd0, 24'd0, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[41] =  { 24'd0, 24'd0, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[42] =  { 24'd0, 24'd0, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd10123859, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[43] =  { 24'd0, 24'd0, 24'd0, 24'd10123859, 24'd10123859, 24'd10123859, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign witch_sprite0[44] =  { 24'd0, 24'd0, 24'd0, 24'd10123859, 24'd10123859, 24'd10123859, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
endmodule // ROM_witch_sprite0