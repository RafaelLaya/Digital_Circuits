/*	ROM module that stores Sprite #3 for dragon
 *		Outputs:
 *			dragon_sprite3			- sprite #3 for dragon
 *
 * Position [x][y][{r,g,b}] contains pixel at (x, y) where r, g, b are 8 bits each
 * (0, 0) is at the top-left
 * Width 45, Height 36, Color-depth 24
*/
module ROM_dragon_sprite3(dragon_sprite3);
	output logic [35:0][23:0] dragon_sprite3 [44:0];
		
	assign dragon_sprite3[0] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[1] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[2] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd16711680, 24'd16711680, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[3] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd16711680, 24'd16711680, 24'd13107200, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[4] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd5046016, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[5] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd13107200, 24'd13107200, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[6] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd13107200, 24'd13107200, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[7] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[8] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[9] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd13107200, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[10] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd16711680, 24'd16711680, 24'd13107200, 24'd13107200, 24'd0, 24'd13107200, 24'd13107200, 24'd13107200, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[11] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd13107200, 24'd16711680, 24'd13107200, 24'd13107200, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[12] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd0, 24'd0, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[13] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd13107200, 24'd13107200, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[14] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[15] =  { 24'd0, 24'd13107200, 24'd13107200, 24'd13107200, 24'd13107200, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[16] =  { 24'd0, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd13107200, 24'd13107200, 24'd13107200, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[17] =  { 24'd0, 24'd0, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[18] =  { 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[19] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[20] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[21] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[22] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[23] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[24] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[25] =  { 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd13107200, 24'd0, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[26] =  { 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd16711680, 24'd13107200, 24'd13107200, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[27] =  { 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd13107200, 24'd13107200, 24'd13107200, 24'd13107200, 24'd13107200, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[28] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[29] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd16711680, 24'd16711680, 24'd16711680, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[30] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd16711680, 24'd16711680, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[31] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd16711680, 24'd16711680, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[32] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd16711680, 24'd13107200, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[33] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd16711680, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[34] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd16711680, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[35] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd16711680, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[36] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[37] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[38] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[39] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[40] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[41] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd13107200, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[42] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[43] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dragon_sprite3[44] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };

endmodule // ROM_dragon_sprite3