/*	ROM module that stores Sprite #0 for dyno in running position
 *		Outputs:
 *			dyno_running_sprite0			- sprite #0 for dyno in running position
 *
 * Position [x][y][{r,g,b}] contains pixel at (x, y) where r, g, b are 8 bits each
 * (0, 0) is at the top-left
 * Width 32, Height 32, Color-depth 24
*/
module ROM_dyno_running_sprite0(dyno_running_sprite0);
	
	output logic [31:0][23:0] dyno_running_sprite0 [0:31];	

	assign dyno_running_sprite0[0] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_running_sprite0[1] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_running_sprite0[2] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_running_sprite0[3] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd0 };
	assign dyno_running_sprite0[4] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd0 };
	assign dyno_running_sprite0[5] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd0 };
	assign dyno_running_sprite0[6] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680 };
	assign dyno_running_sprite0[7] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680 };
	assign dyno_running_sprite0[8] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16711680, 24'd16711680 };
	assign dyno_running_sprite0[9] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite0[10] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite0[11] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd8323072, 24'd8323072, 24'd8323072, 24'd8323072, 24'd16757375, 24'd5011456, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite0[12] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd8323072, 24'd8323072, 24'd8323072, 24'd8323072, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite0[13] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd8323072, 24'd8323072, 24'd0, 24'd0, 24'd0, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd10526880, 24'd10526880, 24'd10526880, 24'd5011456, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite0[14] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd8323072, 24'd8323072, 24'd0, 24'd0, 24'd0, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite0[15] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd8323072, 24'd8323072, 24'd0, 24'd0, 24'd0, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite0[16] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite0[17] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite0[18] =  { 24'd8323072, 24'd8323072, 24'd8323072, 24'd8323072, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd16757375, 24'd16757375, 24'd16711680, 24'd16711680, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite0[19] =  { 24'd8323072, 24'd8323072, 24'd8323072, 24'd8323072, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd16757375, 24'd16757375, 24'd16711680, 24'd16711680, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd16757375, 24'd5011456, 24'd5011456, 24'd5011456 };
	assign dyno_running_sprite0[20] =  { 24'd8323072, 24'd8323072, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16757375, 24'd16757375, 24'd38143, 24'd38143, 24'd16757375, 24'd5011456, 24'd0, 24'd0 };
	assign dyno_running_sprite0[21] =  { 24'd8323072, 24'd8323072, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd5011456, 24'd0, 24'd0, 24'd16711680, 24'd16711680, 24'd16757375, 24'd16757375, 24'd38143, 24'd38143, 24'd16757375, 24'd5011456, 24'd0, 24'd0 };
	assign dyno_running_sprite0[22] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16757375, 24'd16757375, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_running_sprite0[23] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16757375, 24'd16757375, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_running_sprite0[24] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16757375, 24'd16757375, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_running_sprite0[25] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16757375, 24'd16757375, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_running_sprite0[26] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16757375, 24'd16757375, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_running_sprite0[27] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd16711680, 24'd16711680, 24'd0, 24'd0 };
	assign dyno_running_sprite0[28] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd10526880, 24'd16711680, 24'd16711680, 24'd16711680, 24'd16711680, 24'd0, 24'd0 };
	assign dyno_running_sprite0[29] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_running_sprite0[30] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign dyno_running_sprite0[31] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd16766976, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };

endmodule // ROM_dyno_running_sprite0