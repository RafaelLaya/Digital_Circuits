/*	ROM module that stores Sprite for rocket
 *		Outputs:
 *			rocket_sprite		- Sprite for rocket
 *
 * Position [x][y][{r,g,b}] contains pixel at (x, y) where r, g, b are 8 bits each
 * (0, 0) is at the top-left
 * Width 45, Height 36, Color-depth 24
*/
module ROM_rocket_sprite(rocket_sprite);

	output logic [35:0][23:0] rocket_sprite [44:0];

	assign rocket_sprite[0] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[1] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[2] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[3] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[4] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[5] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[6] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[7] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd9571595, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[8] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[9] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[10] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[11] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[12] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[13] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[14] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[15] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[16] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[17] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[18] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[19] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[20] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[21] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[22] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[23] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[24] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[25] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[26] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[27] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[28] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[29] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[30] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[31] =  { 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[32] =  { 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign rocket_sprite[33] =  { 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051 };
	assign rocket_sprite[34] =  { 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051 };
	assign rocket_sprite[35] =  { 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051, 24'd9212051 };

endmodule // ROM_rocket_sprite