/*	ROM module that stores Sprite for eye
 *		Outputs:
 *			eye_sprite			- Sprite for eye
 *
 * Position [x][y][{r,g,b}] contains pixel at (x, y) where r, g, b are 8 bits each
 * (0, 0) is at the top-left
 * Width 45, Height 36, Color-depth 24
*/

module ROM_eye_sprite(eye_sprite);

	output logic [35:0][23:0] eye_sprite [44:0];
		
	assign eye_sprite[0] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[1] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd1315860, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd921102, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[2] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd789516, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[3] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[4] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[5] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[6] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[7] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[8] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[9] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[10] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[11] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[12] =  { 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12191495, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[13] =  { 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd460551, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[14] =  { 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[15] =  { 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[16] =  { 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd3083014, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[17] =  { 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd1973790, 24'd1973790, 24'd1973790, 24'd16740643, 24'd16740643, 24'd16740643, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[18] =  { 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd16740643, 24'd16740643, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd16740643, 24'd16740643, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[19] =  { 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd16740643, 24'd16740643, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd16740643, 24'd16740643, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[20] =  { 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12191495, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd16740643, 24'd16740643, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd16711422, 24'd16711422, 24'd16711422, 24'd1973790, 24'd16740643, 24'd16740643, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[21] =  { 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd16740643, 24'd16740643, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd16711422, 24'd16711422, 24'd16711422, 24'd1973790, 24'd16740643, 24'd16740643, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[22] =  { 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd16740643, 24'd16740643, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd16711422, 24'd16711422, 24'd16711422, 24'd1973790, 24'd16740643, 24'd16740643, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[23] =  { 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd16740643, 24'd16740643, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd16711422, 24'd16711422, 24'd1973790, 24'd1973790, 24'd16740643, 24'd16740643, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[24] =  { 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd16740643, 24'd16740643, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd16740643, 24'd16740643, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd0, 24'd0 };
	assign eye_sprite[25] =  { 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd16740643, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd0, 24'd0 };
	assign eye_sprite[26] =  { 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd16740643, 24'd16740643, 24'd1973790, 24'd1973790, 24'd1973790, 24'd1973790, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd0, 24'd0 };
	assign eye_sprite[27] =  { 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd2887435, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd0, 24'd0 };
	assign eye_sprite[28] =  { 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd0, 24'd0 };
	assign eye_sprite[29] =  { 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd16740643, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[30] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12060423, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd11012359, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[31] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd921102, 24'd12322567, 24'd12322567, 24'd12322567, 24'd789516, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[32] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd0, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[33] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[34] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[35] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[36] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[37] =  { 24'd0, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[38] =  { 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[39] =  { 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[40] =  { 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[41] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[42] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[43] =  { 24'd0, 24'd0, 24'd0, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd12322567, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };
	assign eye_sprite[44] =  { 24'd0, 24'd0, 24'd0, 24'd0, 24'd789516, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0, 24'd0 };

endmodule // eye_sprite